library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library components



entity tb_Bin_BCD is
end;


architecture tb of tb_Bin_BCD is
begin
    stuff!   

